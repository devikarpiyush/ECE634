
  typedef enum bit [1:0] {CSR='b00, DPR='b01, CMDR='b10, FSMR='b11} reg_type_t;

  typedef enum bit {WB_READ_ENB='b0, WB_WRITE_ENB='b1} we_type_t;


